CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 32 408 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 PR
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44679 0
0
13 Logic Switch~
5 24 653 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 CL
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44679 1
0
13 Logic Switch~
5 30 460 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
7 Switch3
-23 -25 26 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44679 2
0
13 Logic Switch~
5 825 673 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
7 Switch4
-23 -26 26 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
44679 3
0
13 Logic Switch~
5 767 308 0 1 11
0 16
0
0 0 21344 0
2 0V
-6 -16 8 -8
7 Switch2
-23 -25 26 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.90029e-315 0
0
13 Logic Switch~
5 25 313 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 CL
-7 -25 7 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90029e-315 5.26354e-315
0
13 Logic Switch~
5 29 48 0 10 11
0 40 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 PR
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90029e-315 5.30499e-315
0
13 Logic Switch~
5 28 166 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
7 Switch1
-23 -25 26 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.90029e-315 5.32571e-315
0
9 Inverter~
13 878 632 0 2 22
0 7 8
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U18A
-36 -4 -8 4
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
4747 0 0
2
5.90029e-315 0
0
9 2-In AND~
219 247 481 0 3 22
0 11 3 10
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U16D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
972 0 0
2
44679 4
0
9 2-In AND~
219 460 497 0 3 22
0 3 4 9
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
3472 0 0
2
44679 5
0
6 74112~
219 133 566 0 7 32
0 13 15 2 15 14 41 3
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U8B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
9998 0 0
2
44679 6
0
6 74112~
219 369 567 0 7 32
0 13 10 2 3 14 42 4
0
0 0 4704 0
5 74112
4 -60 39 -52
4 U10A
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 6 0
1 U
3536 0 0
2
44679 7
0
6 74112~
219 572 566 0 7 32
0 13 9 2 9 14 43 5
0
0 0 4704 0
5 74112
4 -60 39 -52
4 U10B
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 6 0
1 U
4597 0 0
2
44679 8
0
6 74112~
219 733 565 0 7 32
0 13 12 2 3 14 11 6
0
0 0 4704 0
5 74112
4 -60 39 -52
4 U11A
-33 -60 -5 -52
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 7 0
1 U
3835 0 0
2
44679 9
0
7 Pulser~
4 32 539 0 10 12
0 44 45 46 2 0 0 5 5 1
7
0
0 0 4640 0
0
6 Pulser
-20 -28 22 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3670 0 0
2
44679 10
0
9 2-In AND~
219 656 493 0 3 22
0 5 9 12
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U12D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
5616 0 0
2
44679 11
0
9 Inverter~
13 829 268 0 2 22
0 16 17
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U18B
-33 -3 -5 5
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
9323 0 0
2
5.90029e-315 5.34643e-315
0
9 CC 7-Seg~
183 1192 94 0 18 19
10 28 27 26 25 24 23 22 47 48
1 1 0 1 1 0 1 2 2
0
0 0 21104 0
7 AMBERCC
9 -41 58 -33
7 UNIDADE
30 -4 79 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
317 0 0
2
5.90029e-315 5.3568e-315
0
4 4543
219 953 547 0 20 29
0 6 5 4 3 8 7 7 22 23
24 25 26 27 28 0 0 0 0 0
2
0
0 0 4832 0
4 4543
-14 -60 14 -52
3 U13
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 2 3 5 1 7 6 14 15
13 12 11 10 9 4 2 3 5 1
7 6 14 15 13 12 11 10 9 0
65 0 0 0 1 0 0 0
1 U
3108 0 0
2
5.90029e-315 5.36716e-315
0
6 74112~
219 139 202 0 7 32
0 40 20 6 20 21 49 18
0
0 0 4704 0
5 74112
4 -60 39 -52
4 U11B
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 7 0
1 U
4299 0 0
2
5.90029e-315 5.37752e-315
0
6 74112~
219 393 199 0 7 32
0 40 38 6 18 21 50 19
0
0 0 4704 0
5 74112
4 -60 39 -52
4 U15A
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 10 0
1 U
9672 0 0
2
5.90029e-315 5.38788e-315
0
6 74112~
219 647 201 0 7 32
0 40 39 6 18 21 37 29
0
0 0 4704 0
5 74112
4 -60 39 -52
4 U15B
19 -61 47 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 10 0
1 U
7876 0 0
2
5.90029e-315 5.39306e-315
0
9 2-In AND~
219 547 98 0 3 22
0 18 19 39
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
6369 0 0
2
5.90029e-315 5.39824e-315
0
9 2-In AND~
219 291 128 0 3 22
0 37 18 38
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
9172 0 0
2
5.90029e-315 5.40342e-315
0
4 4543
219 900 188 0 14 29
0 51 29 19 18 17 16 16 36 35
34 33 32 31 30
0
0 0 4832 0
4 4543
-14 -60 14 -52
3 U17
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 2 3 5 1 7 6 14 15
13 12 11 10 9 4 2 3 5 1
7 6 14 15 13 12 11 10 9 0
65 0 0 512 1 0 0 0
1 U
7100 0 0
2
5.90029e-315 5.4086e-315
0
9 CC 7-Seg~
183 1096 94 0 18 19
10 30 31 32 33 34 35 36 52 53
1 1 1 1 1 1 0 2 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
6 DEZENA
27 -4 69 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3820 0 0
2
5.90029e-315 5.41378e-315
0
75
3 0 2 0 0 4096 0 14 0 0 18 2
542 539
542 594
3 0 2 0 0 0 0 13 0 0 18 2
339 540
339 594
4 0 3 0 0 12288 0 20 0 0 15 4
921 538
808 538
808 581
690 581
3 7 4 0 0 12416 0 20 13 0 0 6
921 529
793 529
793 571
436 571
436 531
393 531
2 7 5 0 0 4224 0 20 14 0 0 6
921 520
767 520
767 497
681 497
681 530
596 530
3 0 6 0 0 4096 0 23 0 0 8 2
617 174
617 347
3 0 6 0 0 4096 0 22 0 0 8 2
363 172
363 347
0 3 6 0 0 8320 0 0 21 9 0 4
819 511
819 347
109 347
109 175
7 1 6 0 0 0 0 15 20 0 0 3
757 529
757 511
921 511
6 0 7 0 0 8320 0 20 0 0 11 3
921 556
903 556
903 673
7 1 7 0 0 0 0 20 4 0 0 3
921 565
921 673
837 673
1 0 7 0 0 0 0 9 0 0 11 2
881 650
881 673
5 2 8 0 0 8320 0 20 9 0 0 3
921 547
881 547
881 614
4 0 3 0 0 4096 0 13 0 0 15 2
345 549
200 549
4 0 3 0 0 12416 0 15 0 0 21 5
709 547
690 547
690 582
200 582
200 521
2 0 9 0 0 4096 0 14 0 0 17 2
548 530
518 530
0 4 9 0 0 4096 0 0 14 19 0 3
518 497
518 548
548 548
3 0 2 0 0 8320 0 15 0 0 27 4
703 538
703 594
79 594
79 539
3 2 9 0 0 4224 0 11 17 0 0 3
481 497
632 497
632 502
2 3 10 0 0 4224 0 13 10 0 0 3
345 531
245 531
245 504
2 0 3 0 0 0 0 10 0 0 24 3
236 459
200 459
200 521
1 6 11 0 0 8320 0 10 15 0 0 5
254 459
254 458
771 458
771 547
763 547
2 7 4 0 0 0 0 11 13 0 0 3
436 506
436 531
393 531
7 1 3 0 0 0 0 12 11 0 0 5
157 530
157 521
295 521
295 488
436 488
3 2 12 0 0 8320 0 17 15 0 0 4
677 493
695 493
695 529
709 529
1 7 5 0 0 0 0 17 14 0 0 4
632 484
610 484
610 530
596 530
3 4 2 0 0 0 0 12 16 0 0 2
103 539
62 539
1 0 13 0 0 4096 0 12 0 0 31 2
133 503
133 408
1 0 13 0 0 4096 0 13 0 0 31 2
369 504
369 408
1 0 13 0 0 0 0 14 0 0 31 2
572 503
572 408
1 1 13 0 0 4224 0 1 15 0 0 3
44 408
733 408
733 502
5 0 14 0 0 4096 0 12 0 0 35 2
133 578
133 653
5 0 14 0 0 0 0 13 0 0 35 2
369 579
369 653
5 0 14 0 0 0 0 14 0 0 35 2
572 578
572 653
1 5 14 0 0 4224 0 2 15 0 0 3
36 653
733 653
733 577
2 4 15 0 0 8192 0 12 12 0 0 4
109 530
99 530
99 548
109 548
1 2 15 0 0 8320 0 3 12 0 0 4
42 460
99 460
99 530
109 530
0 5 8 0 0 0 0 0 20 0 0 4
922 547
923 547
923 547
921 547
1 0 16 0 0 4096 0 18 0 0 42 2
832 286
832 308
5 2 17 0 0 8320 0 26 18 0 0 3
868 188
832 188
832 250
6 0 16 0 0 8320 0 26 0 0 42 3
868 197
850 197
850 308
1 7 16 0 0 0 0 5 26 0 0 4
779 308
860 308
860 206
868 206
7 4 18 0 0 12416 0 21 26 0 0 6
163 166
221 166
221 243
785 243
785 179
868 179
4 0 18 0 0 0 0 22 0 0 46 2
369 181
178 181
2 7 18 0 0 0 0 25 21 0 0 4
267 137
221 137
221 166
163 166
4 7 18 0 0 0 0 23 21 0 0 5
623 183
623 220
178 220
178 166
163 166
3 7 19 0 0 12416 0 26 22 0 0 6
868 170
730 170
730 133
539 133
539 163
417 163
4 0 20 0 0 4096 0 21 0 0 49 3
115 184
95 184
95 166
1 2 20 0 0 4224 0 8 21 0 0 4
40 166
116 166
116 166
115 166
5 0 21 0 0 4096 0 21 0 0 52 2
139 214
139 313
5 0 21 0 0 4096 0 22 0 0 52 2
393 211
393 313
1 5 21 0 0 4224 0 6 23 0 0 3
37 313
647 313
647 213
8 7 22 0 0 8320 0 20 19 0 0 3
985 565
1207 565
1207 130
9 6 23 0 0 8320 0 20 19 0 0 3
985 556
1201 556
1201 130
10 5 24 0 0 8320 0 20 19 0 0 3
985 547
1195 547
1195 130
11 4 25 0 0 8320 0 20 19 0 0 3
985 538
1189 538
1189 130
12 3 26 0 0 8320 0 20 19 0 0 3
985 529
1183 529
1183 130
13 2 27 0 0 8320 0 20 19 0 0 3
985 520
1177 520
1177 130
14 1 28 0 0 8320 0 20 19 0 0 3
985 511
1171 511
1171 130
7 2 29 0 0 4224 0 23 26 0 0 3
671 165
868 165
868 161
1 14 30 0 0 8320 0 27 26 0 0 3
1075 130
1075 152
932 152
2 13 31 0 0 8320 0 27 26 0 0 3
1081 130
1081 161
932 161
3 12 32 0 0 8320 0 27 26 0 0 3
1087 130
1087 170
932 170
4 11 33 0 0 8320 0 27 26 0 0 3
1093 130
1093 179
932 179
5 10 34 0 0 8320 0 27 26 0 0 3
1099 130
1099 188
932 188
6 9 35 0 0 8320 0 27 26 0 0 3
1105 130
1105 197
932 197
7 8 36 0 0 8320 0 27 26 0 0 3
1111 130
1111 206
932 206
6 1 37 0 0 12416 0 23 25 0 0 6
677 183
681 183
681 68
259 68
259 119
267 119
3 2 38 0 0 4224 0 25 22 0 0 4
312 128
355 128
355 163
369 163
2 3 39 0 0 8320 0 23 24 0 0 4
623 165
608 165
608 98
568 98
7 2 19 0 0 0 0 22 24 0 0 5
417 163
422 163
422 106
523 106
523 107
7 1 18 0 0 0 0 21 24 0 0 4
163 166
178 166
178 89
523 89
1 0 40 0 0 4096 0 21 0 0 75 2
139 139
139 48
1 0 40 0 0 0 0 22 0 0 75 2
393 136
393 48
1 1 40 0 0 4224 0 7 23 0 0 3
41 48
647 48
647 138
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
