CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
54
13 Logic Switch~
5 28 517 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
6 Enable
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3723 0 0
2
44680.5 0
0
13 Logic Switch~
5 59 936 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 OE
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6244 0 0
2
44680.5 0
0
13 Logic Switch~
5 61 855 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 RD
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6421 0 0
2
44680.5 1
0
13 Logic Switch~
5 63 811 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 CS
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7743 0 0
2
44680.5 2
0
13 Logic Switch~
5 29 456 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9840 0 0
2
5.90029e-315 0
0
13 Logic Switch~
5 32 405 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -13 7 -5
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6910 0 0
2
5.90029e-315 5.26354e-315
0
13 Logic Switch~
5 436 69 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 I0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
449 0 0
2
5.90029e-315 5.30499e-315
0
13 Logic Switch~
5 609 76 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 I1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8761 0 0
2
5.90029e-315 5.32571e-315
0
13 Logic Switch~
5 755 82 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 I2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6748 0 0
2
5.90029e-315 5.34643e-315
0
4 4555
219 161 452 0 7 32
0 4 3 2 24 25 26 27
0
0 0 4848 0
4 4555
-14 -60 14 -52
4 U19A
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
65 %D [%16bi %8bi %1i %2i %3i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 3 2 1 4 5 6 7 3 2
1 4 5 6 7 13 14 15 12 11
10 9 0 0 0 0 0 0 0 0
0 19 0
65 0 0 0 2 1 12 0
1 U
7393 0 0
2
44680.5 0
0
9 2-In AND~
219 746 867 0 3 22
0 14 13 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
7699 0 0
2
5.90029e-315 5.3568e-315
0
9 2-In AND~
219 952 882 0 3 22
0 15 13 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
6638 0 0
2
5.90029e-315 5.36716e-315
0
9 2-In AND~
219 606 880 0 3 22
0 11 13 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
4595 0 0
2
5.90029e-315 5.37752e-315
0
12 D Flip-Flop~
219 803 321 0 4 9
0 8 17 52 50
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U24
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9395 0 0
2
5.90029e-315 5.38788e-315
0
12 D Flip-Flop~
219 800 153 0 4 9
0 53 18 54 16
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U5
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3303 0 0
2
5.90029e-315 5.39306e-315
0
12 D Flip-Flop~
219 801 474 0 4 9
0 8 19 55 49
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U4
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4498 0 0
2
5.90029e-315 5.39824e-315
0
12 D Flip-Flop~
219 807 615 0 4 9
0 8 21 56 20
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U2
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9728 0 0
2
5.90029e-315 5.40342e-315
0
12 D Flip-Flop~
219 660 472 0 4 9
0 9 19 57 22
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3789 0 0
2
5.90029e-315 5.4086e-315
0
12 D Flip-Flop~
219 658 320 0 4 9
0 9 17 58 36
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U23
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3978 0 0
2
5.90029e-315 5.41378e-315
0
12 D Flip-Flop~
219 648 617 0 4 9
0 9 21 59 23
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U6
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3494 0 0
2
5.90029e-315 5.41896e-315
0
12 D Flip-Flop~
219 658 153 0 4 9
0 9 18 60 37
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U1
-8 -55 6 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3507 0 0
2
5.90029e-315 5.42414e-315
0
12 D Flip-Flop~
219 486 618 0 4 9
0 10 21 61 12
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U22
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5151 0 0
2
5.90029e-315 5.42933e-315
0
12 D Flip-Flop~
219 491 471 0 4 9
0 10 19 62 40
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U21
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3701 0 0
2
5.90029e-315 5.43192e-315
0
12 D Flip-Flop~
219 491 320 0 4 9
0 10 17 63 46
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U13
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8585 0 0
2
5.90029e-315 5.43451e-315
0
12 D Flip-Flop~
219 491 153 0 4 9
0 10 18 64 47
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U12
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8809 0 0
2
5.90029e-315 5.4371e-315
0
14 Logic Display~
6 359 188 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5993 0 0
2
44680.5 3
0
14 Logic Display~
6 358 363 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8654 0 0
2
44680.5 4
0
14 Logic Display~
6 359 515 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7223 0 0
2
44680.5 5
0
14 Logic Display~
6 364 658 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
44680.5 6
0
14 Logic Display~
6 879 968 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 D0
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3104 0 0
2
44680.5 7
0
14 Logic Display~
6 921 969 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 D1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3296 0 0
2
44680.5 8
0
14 Logic Display~
6 974 972 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 D2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
44680.5 9
0
9 2-In AND~
219 870 698 0 3 22
0 20 27 43
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U18A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
949 0 0
2
44680.5 10
0
9 2-In AND~
219 675 707 0 3 22
0 23 27 32
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U16D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
3371 0 0
2
44680.5 11
0
9 2-In AND~
219 519 706 0 3 22
0 12 27 38
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U16C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
7311 0 0
2
44680.5 12
0
8 4-In OR~
219 924 791 0 5 22
0 48 45 44 43 15
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U17A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 17 0
1 U
3409 0 0
2
44680.5 13
0
8 4-In OR~
219 710 792 0 5 22
0 35 34 33 32 14
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U11B
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 11 0
1 U
3526 0 0
2
44680.5 14
0
8 4-In OR~
219 555 787 0 5 22
0 42 41 39 38 11
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U11A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 11 0
1 U
4129 0 0
2
44680.5 15
0
9 2-In AND~
219 693 561 0 3 22
0 22 26 33
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U16B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
6278 0 0
2
5.90029e-315 5.43969e-315
0
9 2-In AND~
219 907 554 0 3 22
0 49 26 44
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U16A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
3482 0 0
2
5.90029e-315 5.44228e-315
0
9 2-In AND~
219 710 414 0 3 22
0 36 25 34
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U15D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
8323 0 0
2
5.90029e-315 5.44487e-315
0
9 2-In AND~
219 924 413 0 3 22
0 50 25 45
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U15C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
3984 0 0
2
5.90029e-315 5.44746e-315
0
9 2-In AND~
219 539 560 0 3 22
0 40 26 39
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U15B
43 -33 71 -25
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
7622 0 0
2
5.90029e-315 5.45005e-315
0
9 2-In AND~
219 556 410 0 3 22
0 46 25 41
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U15A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
816 0 0
2
5.90029e-315 5.45264e-315
0
9 2-In AND~
219 942 241 0 3 22
0 16 24 48
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
4656 0 0
2
5.90029e-315 5.45523e-315
0
9 2-In AND~
219 727 239 0 3 22
0 37 24 35
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
6356 0 0
2
5.90029e-315 5.45782e-315
0
9 2-In AND~
219 570 238 0 3 22
0 47 24 42
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
7479 0 0
2
5.90029e-315 5.46041e-315
0
9 2-In AND~
219 397 647 0 3 22
0 51 27 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
5690 0 0
2
5.90029e-315 5.463e-315
0
9 2-In AND~
219 389 491 0 3 22
0 51 26 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
5617 0 0
2
5.90029e-315 5.46559e-315
0
9 2-In AND~
219 387 351 0 3 22
0 51 25 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3903 0 0
2
5.90029e-315 5.46818e-315
0
9 2-In AND~
219 391 162 0 3 22
0 51 24 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
4452 0 0
2
5.90029e-315 5.47077e-315
0
5 7415~
219 477 927 0 4 22
0 29 28 30 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 10 0
1 U
6282 0 0
2
5.90029e-315 5.47207e-315
0
9 2-In AND~
219 353 759 0 3 22
0 28 31 51
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U9A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
7187 0 0
2
5.90029e-315 5.48372e-315
0
5 4069~
219 358 829 0 2 22
0 29 31
0
0 0 624 90
4 4069
-7 -24 21 -16
3 U8E
16 -2 37 6
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 8 0
1 U
6866 0 0
2
5.90029e-315 5.48502e-315
0
92
3 1 2 0 0 8336 0 10 1 0 0 4
123 452
72 452
72 517
40 517
1 2 3 0 0 12416 0 5 10 0 0 4
41 456
58 456
58 434
129 434
1 1 4 0 0 12416 0 6 10 0 0 4
44 405
58 405
58 425
129 425
3 1 5 0 0 8320 0 12 32 0 0 3
973 882
974 882
974 958
3 1 6 0 0 8320 0 11 31 0 0 4
767 867
767 892
921 892
921 955
3 1 7 0 0 8320 0 13 30 0 0 4
627 880
627 906
879 906
879 954
1 0 8 0 0 4096 0 14 0 0 9 2
779 285
756 285
1 0 8 0 0 0 0 16 0 0 9 2
777 438
756 438
1 1 8 0 0 8320 0 9 17 0 0 4
755 94
756 94
756 579
783 579
1 0 9 0 0 4096 0 18 0 0 42 2
636 436
608 436
1 0 9 0 0 0 0 19 0 0 42 2
634 284
608 284
1 0 9 0 0 0 0 21 0 0 42 2
634 117
608 117
1 0 10 0 0 4096 0 25 0 0 40 2
467 117
435 117
1 0 10 0 0 0 0 24 0 0 40 2
467 284
435 284
1 0 10 0 0 0 0 23 0 0 40 2
467 435
435 435
5 1 11 0 0 4224 0 38 13 0 0 3
558 817
558 871
582 871
4 1 12 0 0 8320 0 22 35 0 0 3
510 582
526 582
526 684
2 0 13 0 0 4096 0 13 0 0 20 2
582 889
582 927
2 0 13 0 0 4096 0 11 0 0 20 2
722 876
722 927
4 2 13 0 0 4224 0 52 12 0 0 3
498 927
928 927
928 891
5 1 14 0 0 4224 0 37 11 0 0 3
713 822
713 858
722 858
5 1 15 0 0 4224 0 36 12 0 0 3
927 821
927 873
928 873
4 1 16 0 0 4224 0 15 45 0 0 3
824 117
949 117
949 219
2 0 17 0 0 4096 0 19 0 0 26 2
634 302
634 351
2 0 17 0 0 0 0 24 0 0 26 2
467 302
467 351
3 2 17 0 0 4224 0 50 14 0 0 3
408 351
779 351
779 303
2 0 18 0 0 4096 0 21 0 0 29 2
634 135
634 162
2 0 18 0 0 0 0 25 0 0 29 2
467 135
467 162
3 2 18 0 0 4224 0 51 15 0 0 3
412 162
776 162
776 135
2 0 19 0 0 4096 0 23 0 0 32 2
467 453
467 491
2 0 19 0 0 0 0 18 0 0 32 2
636 454
636 491
3 2 19 0 0 4224 0 49 16 0 0 3
410 491
777 491
777 456
4 1 20 0 0 8320 0 17 33 0 0 3
831 579
877 579
877 676
2 0 21 0 0 4096 0 22 0 0 36 2
462 600
462 647
2 0 21 0 0 4096 0 20 0 0 36 2
624 599
624 647
3 2 21 0 0 4224 0 48 17 0 0 3
418 647
783 647
783 597
4 0 22 0 0 0 0 18 0 0 53 2
684 436
684 436
4 1 23 0 0 8320 0 20 34 0 0 3
672 581
682 581
682 685
1 0 9 0 0 0 0 20 0 0 42 2
624 581
624 581
1 1 10 0 0 8320 0 7 22 0 0 6
436 81
435 81
435 440
436 440
436 582
462 582
4 0 12 0 0 0 0 22 0 0 0 2
510 582
516 582
1 0 9 0 0 12416 0 8 0 0 0 5
609 88
609 117
608 117
608 581
630 581
1 0 24 0 0 4096 0 26 0 0 92 2
359 206
359 205
1 0 25 0 0 4096 0 27 0 0 86 2
358 381
358 379
1 0 26 0 0 4096 0 28 0 0 84 2
359 533
359 533
1 0 27 0 0 4096 0 29 0 0 77 2
364 676
364 679
2 0 28 0 0 4096 0 52 0 0 51 3
453 927
296 927
296 811
0 1 29 0 0 8192 0 0 52 50 0 3
360 854
360 918
453 918
1 3 30 0 0 4224 0 2 52 0 0 2
71 936
453 936
1 1 29 0 0 4224 0 3 54 0 0 5
73 855
360 855
360 854
361 854
361 847
1 1 28 0 0 4224 0 4 53 0 0 3
75 811
343 811
343 780
2 2 31 0 0 4224 0 54 53 0 0 2
361 811
361 780
0 1 22 0 0 8320 0 0 39 0 0 3
680 436
700 436
700 539
2 0 27 0 0 4096 0 34 0 0 77 2
664 685
664 679
2 0 26 0 0 4096 0 39 0 0 84 2
682 539
682 533
2 0 25 0 0 4096 0 41 0 0 86 2
699 392
699 379
2 0 24 0 0 4096 0 46 0 0 92 2
716 217
716 205
3 4 32 0 0 4224 0 34 37 0 0 3
673 730
673 772
699 772
3 3 33 0 0 4224 0 39 37 0 0 4
691 584
691 767
708 767
708 772
3 2 34 0 0 4224 0 41 37 0 0 4
708 437
708 763
717 763
717 772
3 1 35 0 0 8320 0 46 37 0 0 3
725 262
726 262
726 772
4 1 36 0 0 8320 0 19 41 0 0 3
682 284
717 284
717 392
4 1 37 0 0 8320 0 21 46 0 0 3
682 117
734 117
734 217
2 0 24 0 0 0 0 47 0 0 92 2
559 216
559 205
2 0 25 0 0 0 0 44 0 0 86 2
545 388
545 379
3 4 38 0 0 4224 0 35 38 0 0 4
517 729
517 760
544 760
544 767
2 0 27 0 0 0 0 35 0 0 77 2
508 684
508 679
3 3 39 0 0 4224 0 43 38 0 0 4
537 583
537 756
553 756
553 767
2 0 26 0 0 0 0 43 0 0 84 2
528 538
528 533
4 1 40 0 0 12416 0 23 43 0 0 4
515 435
515 436
546 436
546 538
3 2 41 0 0 8320 0 44 38 0 0 3
554 433
562 433
562 767
3 1 42 0 0 8320 0 47 38 0 0 3
568 261
571 261
571 767
2 0 27 0 0 4096 0 48 0 0 77 2
373 656
373 679
3 4 43 0 0 4224 0 33 36 0 0 4
868 721
868 768
913 768
913 771
3 3 44 0 0 4224 0 40 36 0 0 4
905 577
905 764
922 764
922 771
3 2 45 0 0 4224 0 42 36 0 0 4
922 436
922 758
931 758
931 771
7 2 27 0 0 12416 0 10 33 0 0 5
193 425
243 425
243 679
859 679
859 676
4 1 46 0 0 8320 0 24 44 0 0 3
515 284
563 284
563 388
4 1 47 0 0 8320 0 25 47 0 0 3
515 117
577 117
577 216
1 3 48 0 0 4224 0 36 45 0 0 2
940 771
940 264
4 1 49 0 0 8320 0 16 40 0 0 3
825 438
914 438
914 532
4 1 50 0 0 8320 0 14 42 0 0 3
827 285
931 285
931 391
2 0 26 0 0 4096 0 49 0 0 84 2
365 500
365 533
6 2 26 0 0 12416 0 10 40 0 0 5
193 434
252 434
252 533
896 533
896 532
2 0 25 0 0 4096 0 50 0 0 86 2
363 360
363 379
5 2 25 0 0 12416 0 10 42 0 0 5
193 443
235 443
235 379
913 379
913 391
1 0 51 0 0 4096 0 48 0 0 90 2
373 638
352 638
1 0 51 0 0 0 0 49 0 0 90 2
365 482
352 482
1 0 51 0 0 0 0 50 0 0 90 2
363 342
352 342
3 1 51 0 0 4224 0 53 51 0 0 3
352 735
352 153
367 153
2 0 24 0 0 4096 0 51 0 0 92 2
367 171
367 205
4 2 24 0 0 12416 0 10 45 0 0 5
193 452
227 452
227 205
931 205
931 219
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
